../../lib/pcores/reconos_fifo_async_v1_00_a/hdl/vhdl/reconos_fifo_async.vhd